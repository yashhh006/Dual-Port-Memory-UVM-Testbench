`include "uvm_pkg.sv"
import uvm_pkg::*;

`include "memory.sv"
`include "mem_comm.sv"
`include "mem_intf.sv"
`include "mem_tx.sv"
`include "mem_tx3.sv"
`include "mem_seq.sv"
`include "mem_sqr.sv"
`include "mem_drv.sv"
`include "mem_cov.sv"
`include "mem_mon.sv"
`include "mem_agent.sv"
`include "mem_tx2.sv"
`include "mem_seq2.sv"
`include "mem_sqr2.sv"
`include "mem_drv2.sv"
`include "mem_drv3.sv"
`include "mem_cov2.sv"
`include "mem_mon2.sv"
`include "mem_agent2.sv"
`include "mem_sbd.sv"
`include "mem_env.sv"
`include "mem_test.sv"

`include "top.sv"