//Two always block for two ports

//Flag mechanism to prevent both ports trying ot access the same location

//bit [width-1:0]flag[depth-1:0];