`include "list.svh"